//------------------------------------------------------------------------------
// Copyright (c) 2021 by Ando Ki.
// All rights reserved by Ando Ki.
//------------------------------------------------------------------------------
// cosim_bfm_axi_dpi.sv
//------------------------------------------------------------------------------

`define COSIM_DPI
`undef  COSIM_VPI
`include "cosim_bfm_axi_core.v"

//------------------------------------------------------------------------------
// Revision history
//
// 2021.07.01: Started by Ando Ki (andoki@gmail.com)
//------------------------------------------------------------------------------
